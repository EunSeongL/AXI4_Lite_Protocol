`timescale 1ns / 1ps

module AXI4_Lite_Master (
    // global signals
    input logic ACLK,
    input logic ARESETn,
    // Write Transfer, AW Channel
    output logic [3:0] AWADDR,
    output logic       AWVALID,
    input  logic       AWREADY,
    // Write Transfer, W Channel
    output logic [31:0] WDATA,
    output logic        WVALID,
    input logic         WREADY,
    // Write Transfer, B Channel
    input logic [1:0] BRESP,
    input logic       BVALID,
    output logic      BREADY,
    // READ Transfer, AR Channel
    output logic [3:0] ARADDR,
    output logic       ARVALID,
    input logic        ARREADY,
    // READ Transfer, R Channel
    input logic  [31:0] RDATA,
    input logic  [1:0] RRESP,
    input logic         RVALID,
    output logic        RREADY,
    // internal signals
    input logic [3:0] addr,
    input logic       write,
    input logic [31:0] wdata,
    output logic [31:0] rdata,
    input logic transfer,
    output logic ready
);

    // Write Transaction, AW (Write Addr)channel Transfer
    typedef enum {
        AW_IDLE,
        AW_VALID
    } aw_state_e;
    
    aw_state_e aw_state, aw_state_next;
    logic [3:0] temp_awaddr_reg, temp_awaddr_next;

    always_ff @(posedge ACLK or posedge ARESETn) begin
        if(!ARESETn) begin
            AW_IDLE <= aw_state;
            temp_awaddr_reg <= 0;
        end
        else begin
            aw_state <= aw_state_next;
            temp_awaddr_reg <= temp_awaddr_next;
        end
    end

    always_comb begin
        aw_state_next = aw_state;
        AWADDR = temp_awaddr_reg;
        AWVALID = 1'b0;
        case (aw_state)
            AW_IDLE: begin
                AWVALID = 0;
                temp_wdata_next = addr;
                if(transfer & write) begin
                    aw_state_next = AW_VALID;
                end
            end
            AW_VALID: begin
                AWVALID = 1'b1;
                AWADDR = temp_awaddr_reg;
                if(AWREADY) begin
                    aw_state_next = AW_IDLE;
                end
            end
        endcase
    end
    // Write Transaction, W (Write Data) Channel Transfer
    typedef enum {
        W_IDLE,
        W_VALID
    } w_state_e;
    
    w_state_e w_state, w_state_next;
    logic [31:0] temp_wdata_next, temp_wdata_reg;

    always_ff @(posedge ACLK or posedge ARESETn) begin
        if(!ARESETn) begin
            W_IDLE <= w_state;
            temp_wdata_reg <= 0;
        end
        else begin
            w_state <= w_state_next;
            temp_wdata_reg <= temp_wdata_next;
        end
    end

    always_comb begin
        w_state_next = w_state;
        WDATA = temp_wdata_reg;
        WVALID = 1'b0;
        case (w_state)
            W_IDLE: begin
                WVALID = 0;
                temp_wdata_next = wdata;
                if(transfer & write) begin
                    w_state_next = W_VALID;
                end
            end
            W_VALID: begin
                WVALID = 1'b1;
                WDATA = temp_wdata_reg;
                if(WREADY) begin
                    w_state_next = W_IDLE;
                end
            end
        endcase
    end
    // WRITE Transaction, B Channel Transfer BRESP = 2'b00 : OKAY 
    typedef enum {
        B_IDLE,
        B_READY
    } b_state_e;
    
    b_state_e b_state, b_state_next;

    always_ff @(posedge ACLK or posedge ARESETn) begin
        if(!ARESETn) begin
            B_IDLE <= b_state;
        end
        else begin
            b_state <= b_state_next;
        end
    end

    always_comb begin
        b_state_next = b_state;
        BREADY = 1'b0;
        w_ready = 1'b0;
        case (b_state)
            B_IDLE: begin
                if(WVALID) begin
                    BREADY = 1'b0;
                    w_ready = 1'b0;
                    b_state_next = B_READY;
                end
            end
            B_READY: begin
                BREADY = 1'b1;
                if(BVALID) begin
                    w_ready = 1'b1;
                    b_state_next = B_IDLE;
                end
            end
        endcase
    end

    // READ Transaction, AR Channel Transfer
    typedef enum {
        AR_IDLE,
        AR_VALID
    } ar_state_e;

    ar_state_e ar_state, ar_state_next;
    logic [3:0] temp_araddr_reg, temp_araddr_next;

    always_ff @(posedge ACLK or posedge ARESETn) begin 
        if(!ARESET) begin
            ar_state <= AR_IDLE;
            temp_araddr_reg <= 0;
        end
        else begin
            ar_state <= ar_state_next;
            temp_awaddr_reg <= temp_araddr_next;
        end
    end

    always_comb begin
        ar_state_next = ar_state;
        ARADDR = temp_araddr_reg;
        case (ar_state)
            AR_IDLE: begin
                AR_VALID = 1'b0;
                temp_araddr_next = addr;
                if(ready & (!write))begin
                    ar_state_next = AR_VALID;        
                end
            end
            AR_VALID: begin
                AR_VALID = 1'b1;
                ARADDR = temp_araddr_reg;
                if(ARREADY) begin
                    ar_state_next = AR_IDLE;
                end
            end
        endcase
    end

    // READ Transaction, R Channel Transfer
    typedef enum {
        R_IDLE,
        R_READY
    } r_state_e;

    r_state_e r_state, r_state_next;

    always_ff @(posedge ACLK or posedge ARESETn) begin
        if(!ARESETn)begin
            r_state <= R_IDLE;
        end
        else begin
            r_state <= r_state_next;
        end
    end

    always_comb begin
        r_state_next = r_state;
        RREADY = 1'b0;
        r_ready = 1'b0;
        case (r_state)
            R_IDLE:begin
                r_ready = 1'b0;
                RREADY = 1'b0;
                if(ARVALID) r_state_next = R_READY;
            end
            R_READY:begin
                RREADY = 1'b1;
                if(RVALID) begin
                    r_state_next = R_IDLE;
                    r_ready = 1'b1;
                    rdata = RDATA;
                end
            end 
        endcase
    end
endmodule